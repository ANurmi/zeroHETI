module zeroheti_core import zeroheti_pkg::AddrMap; #(
  zeroheti_pkg::core_cfg_t Cfg = zeroheti_pkg::DefaultCfg
)(
  input  logic clk_i,
  input  logic rst_ni,
  input  logic testmode_i,
  input  logic jtag_tck_i,
  input  logic jtag_tms_i,
  input  logic jtag_trst_ni,
  input  logic jtag_td_i,
  output logic jtag_td_o,
  APB.Master   apb_mgr
);

localparam int unsigned NumSbrPorts  = 32'd3;
localparam int unsigned NumMgrPorts  = 32'd5;
localparam int unsigned NumAddrRules = 32'd5;

localparam bit [NumSbrPorts-1:0][NumMgrPorts-1:0] Connectivity = '1; // TODO: minimal required connectivity
/*
obi_cut_intf i_obi_cut (
  .clk_i,
  .rst_ni,
  .obi_s  (sbr_bus[3]),
  .obi_m  (apb_cut)
);*/

obi_to_apb_intf i_obi_to_apb (
  .clk_i,
  .rst_ni,
  .obi_i  (sbr_bus[3]),
  .apb_o  (apb_mgr)
);

typedef struct packed {
  int unsigned idx;
  logic [31:0] start_addr;
  logic [31:0] end_addr;
} addr_map_rule_t;

localparam addr_map_rule_t [NumAddrRules-1:0] CoreAddrMap = '{
  '{idx: 0, start_addr: AddrMap.dbg.base,  end_addr: AddrMap.dbg.last},
  '{idx: 1, start_addr: AddrMap.imem.base, end_addr: AddrMap.imem.last},
  '{idx: 2, start_addr: AddrMap.dmem.base, end_addr: AddrMap.dmem.last},
  // TODO: map other APB peripherals
  '{idx: 3, start_addr: AddrMap.clic.base, end_addr: AddrMap.mtimer.last},
  '{idx: 4, start_addr: AddrMap.ext.base,  end_addr: AddrMap.ext.last}
};

OBI_BUS mgr_bus [NumSbrPorts]();
OBI_BUS sbr_bus [NumMgrPorts]();
//OBI_BUS apb_cut ();

logic debug_req;

obi_xbar_intf #(
  .NumSbrPorts     (NumSbrPorts),
  .NumMgrPorts     (NumMgrPorts),
  .NumMaxTrans     (32'd1),
  .NumAddrRules    (NumAddrRules),
  .addr_map_rule_t (addr_map_rule_t),
  .Connectivity    (Connectivity)
) i_xbar (
  .clk_i,
  .rst_ni,
  .testmode_i,
  .addr_map_i       (CoreAddrMap),
  .en_default_idx_i (3'b0),
  .default_idx_i    (9'b0),
  .sbr_ports        (mgr_bus),
  .mgr_ports        (sbr_bus)
);


`ifndef SYNTHESIS
ibex_top_tracing #(
`else
ibex_top #(
`endif
  .PMPEnable        (0),
  .PMPGranularity   (0),
  .PMPNumRegions    (4),
  .MHPMCounterNum   (0),
  .MHPMCounterWidth (40),
  .RV32E            (Cfg.rve),
  .RV32M            (ibex_pkg::RV32MFast),
  .RV32B            (ibex_pkg::RV32BNone),
  .WritebackStage   (Cfg.wb_stage),
  .RegFile          (ibex_pkg::RegFileWindowFF),
  .ICache           (1'b0),
  .ICacheECC        (1'b0),
  .ICacheScramble   (1'b0),
  .BranchPredictor  (1'b0),
  .SecureIbex       (1'b0),
  .CLIC             (1'b1),
  .HardwareStacking (1'b0),
  .NumInterrupts    (Cfg.num_irqs),
  .RndCnstLfsrSeed  (ibex_pkg::RndCnstLfsrSeedDefault),
  .RndCnstLfsrPerm  (ibex_pkg::RndCnstLfsrPermDefault),
  .DbgTriggerEn     (0),
  .DmHaltAddr       (dm::HaltAddress),
  .DmExceptionAddr  (dm::ExceptionAddress),
  .MClicBaseAddr    (zeroheti_pkg::AddrMap.clic.base),
  .BranchTargetALU  (Cfg.bt_alu)
) i_rt_ibex (
  .clk_i,
  .rst_ni,
  .scan_rst_ni            (1'b0),
  .ram_cfg_i              (10'b0),
  .hart_id_i              (Cfg.hart_id),
  .test_en_i              (testmode_i),
  .boot_addr_i            (Cfg.boot_addr),

  .instr_req_o            (mgr_bus[1].req),
  .instr_addr_o           (mgr_bus[1].addr),
  .instr_gnt_i            (mgr_bus[1].gnt),
  .instr_rvalid_i         (mgr_bus[1].rvalid),
  .instr_rdata_i          (mgr_bus[1].rdata),
  .instr_rdata_intg_i     (7'b0),
  .instr_err_i            (mgr_bus[1].err),

  .data_req_o             (mgr_bus[2].req),
  .data_gnt_i             (mgr_bus[2].gnt),
  .data_rvalid_i          (mgr_bus[2].rvalid),
  .data_we_o              (mgr_bus[2].we),
  .data_be_o              (mgr_bus[2].be),
  .data_addr_o            (mgr_bus[2].addr),
  .data_wdata_o           (mgr_bus[2].wdata),
  .data_rdata_i           (mgr_bus[2].rdata),
  .data_err_i             (mgr_bus[2].err),
  .data_rdata_intg_i      (7'b0),
  .data_wdata_intg_o      (),

  .irq_is_pcs_i           (),
  .irq_i                  (),
  .irq_id_o               (),
  .irq_ack_o              (),
  .irq_level_i            (),
  .irq_shv_i              (),
  .irq_priv_i             (),

  .scramble_key_valid_i   (1'b0),
  .scramble_key_i         (128'b0),
  .scramble_nonce_i       (64'b0),
  .scramble_req_o         (),

  .debug_req_i            (debug_req),
  .debug_mode_o           (),
  .crash_dump_o           (),
  .double_fault_seen_o    (),
  .fetch_enable_i         (4'b0101),
  .core_sleep_o           (),

  .alert_minor_o          (),
  .alert_major_internal_o (),
  .alert_major_bus_o      ()
);

zeroheti_dbg_wrapper #(

) i_debug (
  .clk_i,
  .rst_ni,
  .testmode_i,
  .jtag_tck_i,
  .jtag_tms_i,
  .jtag_trst_ni,
  .jtag_td_i,
  .jtag_td_o,
  .ndmreset_o  (),
  .debug_req_o (debug_req),
  .mem_sbr     (sbr_bus[0]),
  .sba_mgr     (mgr_bus[0])
);

obi_sram_intf #(
  .BaseAddr (AddrMap.imem.base)
) i_imem (
  .clk_i,
  .rst_ni,
  .sbr     (sbr_bus[1])
);

obi_sram_intf #(
  .BaseAddr (AddrMap.dmem.base)
) i_dmem (
  .clk_i,
  .rst_ni,
  .sbr     (sbr_bus[2])
);

endmodule : zeroheti_core

