module zeroheti_dbg_wrapper #()();
endmodule : zeroheti_dbg_wrapper

