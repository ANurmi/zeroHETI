module obi_sram_intf #()(
  input logic clk_i,
  input logic rst_ni
);

/*
obi_sram_shim #(
) i_shim (
  .clk_i,
  .rst_ni,
  .obi_req_i (),
  .obi_rsp_o (),
  .req_o     (),
  .gnt_i     ()
  .we_o      (),
  .addr_o    ()
);*/

endmodule : obi_sram_intf

