module zeroheti_compliance #()();
endmodule : zeroheti_compliance

